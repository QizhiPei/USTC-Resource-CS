
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hb77c7952;
    ram_cell[       1] = 32'h0;  // 32'h996142f5;
    ram_cell[       2] = 32'h0;  // 32'h968cdec9;
    ram_cell[       3] = 32'h0;  // 32'h06e2db2f;
    ram_cell[       4] = 32'h0;  // 32'ha8192a9e;
    ram_cell[       5] = 32'h0;  // 32'h721a6192;
    ram_cell[       6] = 32'h0;  // 32'had036e69;
    ram_cell[       7] = 32'h0;  // 32'h9d42a8f3;
    ram_cell[       8] = 32'h0;  // 32'h1d7b5c10;
    ram_cell[       9] = 32'h0;  // 32'hd2cab7bb;
    ram_cell[      10] = 32'h0;  // 32'h527b2abe;
    ram_cell[      11] = 32'h0;  // 32'hd961cf2c;
    ram_cell[      12] = 32'h0;  // 32'hd73618f5;
    ram_cell[      13] = 32'h0;  // 32'h14dfb33f;
    ram_cell[      14] = 32'h0;  // 32'h17e4b572;
    ram_cell[      15] = 32'h0;  // 32'h8a978fc5;
    ram_cell[      16] = 32'h0;  // 32'h77e5359a;
    ram_cell[      17] = 32'h0;  // 32'h704b342f;
    ram_cell[      18] = 32'h0;  // 32'haac4dd09;
    ram_cell[      19] = 32'h0;  // 32'hd66493aa;
    ram_cell[      20] = 32'h0;  // 32'h5bce4ca4;
    ram_cell[      21] = 32'h0;  // 32'h41048642;
    ram_cell[      22] = 32'h0;  // 32'h7f077004;
    ram_cell[      23] = 32'h0;  // 32'h34862689;
    ram_cell[      24] = 32'h0;  // 32'h30338881;
    ram_cell[      25] = 32'h0;  // 32'hacf19748;
    ram_cell[      26] = 32'h0;  // 32'hd2dc8d86;
    ram_cell[      27] = 32'h0;  // 32'h72c74f3c;
    ram_cell[      28] = 32'h0;  // 32'h486c795c;
    ram_cell[      29] = 32'h0;  // 32'h7296e90a;
    ram_cell[      30] = 32'h0;  // 32'h4ec60e29;
    ram_cell[      31] = 32'h0;  // 32'h906e7624;
    ram_cell[      32] = 32'h0;  // 32'h18469a53;
    ram_cell[      33] = 32'h0;  // 32'h9d7805d4;
    ram_cell[      34] = 32'h0;  // 32'hefb2f25f;
    ram_cell[      35] = 32'h0;  // 32'hc99c01a2;
    ram_cell[      36] = 32'h0;  // 32'h59440d45;
    ram_cell[      37] = 32'h0;  // 32'h3c0af49a;
    ram_cell[      38] = 32'h0;  // 32'h5ae270b3;
    ram_cell[      39] = 32'h0;  // 32'he8e2e4d6;
    ram_cell[      40] = 32'h0;  // 32'hdc58ca7c;
    ram_cell[      41] = 32'h0;  // 32'hbaebddf1;
    ram_cell[      42] = 32'h0;  // 32'h197266f9;
    ram_cell[      43] = 32'h0;  // 32'h0fd97961;
    ram_cell[      44] = 32'h0;  // 32'h3a4449be;
    ram_cell[      45] = 32'h0;  // 32'had04005f;
    ram_cell[      46] = 32'h0;  // 32'h0a129d5c;
    ram_cell[      47] = 32'h0;  // 32'h912461a3;
    ram_cell[      48] = 32'h0;  // 32'h2b7681ce;
    ram_cell[      49] = 32'h0;  // 32'h95dc300f;
    ram_cell[      50] = 32'h0;  // 32'h86fd2aa2;
    ram_cell[      51] = 32'h0;  // 32'hbd828022;
    ram_cell[      52] = 32'h0;  // 32'h7b0f888f;
    ram_cell[      53] = 32'h0;  // 32'h313c12f2;
    ram_cell[      54] = 32'h0;  // 32'ha1cc4472;
    ram_cell[      55] = 32'h0;  // 32'hb3de91b1;
    ram_cell[      56] = 32'h0;  // 32'h4e5c47e2;
    ram_cell[      57] = 32'h0;  // 32'hb2dbac62;
    ram_cell[      58] = 32'h0;  // 32'hcb01db3a;
    ram_cell[      59] = 32'h0;  // 32'h83242af6;
    ram_cell[      60] = 32'h0;  // 32'hff99c846;
    ram_cell[      61] = 32'h0;  // 32'h8555df2b;
    ram_cell[      62] = 32'h0;  // 32'h8af2f0a6;
    ram_cell[      63] = 32'h0;  // 32'h5a1d2f25;
    ram_cell[      64] = 32'h0;  // 32'h923e642b;
    ram_cell[      65] = 32'h0;  // 32'h0bf3c54d;
    ram_cell[      66] = 32'h0;  // 32'h2dbfae38;
    ram_cell[      67] = 32'h0;  // 32'hec9342bc;
    ram_cell[      68] = 32'h0;  // 32'h8890a55a;
    ram_cell[      69] = 32'h0;  // 32'h8db547c8;
    ram_cell[      70] = 32'h0;  // 32'hff27e884;
    ram_cell[      71] = 32'h0;  // 32'h174e2dcd;
    ram_cell[      72] = 32'h0;  // 32'h08ebd670;
    ram_cell[      73] = 32'h0;  // 32'h30c60a98;
    ram_cell[      74] = 32'h0;  // 32'h9e818829;
    ram_cell[      75] = 32'h0;  // 32'h61592ba5;
    ram_cell[      76] = 32'h0;  // 32'h7e29de1b;
    ram_cell[      77] = 32'h0;  // 32'hc7a6d422;
    ram_cell[      78] = 32'h0;  // 32'h7f350774;
    ram_cell[      79] = 32'h0;  // 32'hbc613adc;
    ram_cell[      80] = 32'h0;  // 32'he7ebb109;
    ram_cell[      81] = 32'h0;  // 32'he2c118ff;
    ram_cell[      82] = 32'h0;  // 32'ha43a4b03;
    ram_cell[      83] = 32'h0;  // 32'h6d5a2650;
    ram_cell[      84] = 32'h0;  // 32'h915e8715;
    ram_cell[      85] = 32'h0;  // 32'h8280333a;
    ram_cell[      86] = 32'h0;  // 32'hd7498bf3;
    ram_cell[      87] = 32'h0;  // 32'h87f04e5a;
    ram_cell[      88] = 32'h0;  // 32'h489cd14a;
    ram_cell[      89] = 32'h0;  // 32'h3436725b;
    ram_cell[      90] = 32'h0;  // 32'h6dc9b2a7;
    ram_cell[      91] = 32'h0;  // 32'ha0dfe019;
    ram_cell[      92] = 32'h0;  // 32'hbc102b7c;
    ram_cell[      93] = 32'h0;  // 32'h80b4f812;
    ram_cell[      94] = 32'h0;  // 32'he644fa8f;
    ram_cell[      95] = 32'h0;  // 32'hb18c9f2f;
    ram_cell[      96] = 32'h0;  // 32'h9d041371;
    ram_cell[      97] = 32'h0;  // 32'h904d1c29;
    ram_cell[      98] = 32'h0;  // 32'he6fcd480;
    ram_cell[      99] = 32'h0;  // 32'h263a4a3f;
    ram_cell[     100] = 32'h0;  // 32'h1c76a971;
    ram_cell[     101] = 32'h0;  // 32'h97ba289c;
    ram_cell[     102] = 32'h0;  // 32'hf3caabbe;
    ram_cell[     103] = 32'h0;  // 32'h58b393b7;
    ram_cell[     104] = 32'h0;  // 32'ha9ca3330;
    ram_cell[     105] = 32'h0;  // 32'h4c2fbca5;
    ram_cell[     106] = 32'h0;  // 32'h62fa1887;
    ram_cell[     107] = 32'h0;  // 32'h5af107de;
    ram_cell[     108] = 32'h0;  // 32'hf04401c4;
    ram_cell[     109] = 32'h0;  // 32'h1bad0739;
    ram_cell[     110] = 32'h0;  // 32'h8d729c34;
    ram_cell[     111] = 32'h0;  // 32'h3f32e452;
    ram_cell[     112] = 32'h0;  // 32'h7da94a6d;
    ram_cell[     113] = 32'h0;  // 32'hea274402;
    ram_cell[     114] = 32'h0;  // 32'h7cb88129;
    ram_cell[     115] = 32'h0;  // 32'hcb616742;
    ram_cell[     116] = 32'h0;  // 32'h5824392e;
    ram_cell[     117] = 32'h0;  // 32'h7489ec57;
    ram_cell[     118] = 32'h0;  // 32'hf578f40a;
    ram_cell[     119] = 32'h0;  // 32'heaada014;
    ram_cell[     120] = 32'h0;  // 32'hbd4249a6;
    ram_cell[     121] = 32'h0;  // 32'h3e57608f;
    ram_cell[     122] = 32'h0;  // 32'h4619e2f9;
    ram_cell[     123] = 32'h0;  // 32'h98f51cbe;
    ram_cell[     124] = 32'h0;  // 32'h0219c6bc;
    ram_cell[     125] = 32'h0;  // 32'hc89de25b;
    ram_cell[     126] = 32'h0;  // 32'h33ba5a68;
    ram_cell[     127] = 32'h0;  // 32'heda25518;
    ram_cell[     128] = 32'h0;  // 32'hbea89f51;
    ram_cell[     129] = 32'h0;  // 32'ha002c9b8;
    ram_cell[     130] = 32'h0;  // 32'h6d1e7d2e;
    ram_cell[     131] = 32'h0;  // 32'h3ce3d204;
    ram_cell[     132] = 32'h0;  // 32'h95e35478;
    ram_cell[     133] = 32'h0;  // 32'hd7b97418;
    ram_cell[     134] = 32'h0;  // 32'hb19c3f67;
    ram_cell[     135] = 32'h0;  // 32'hc3d9668c;
    ram_cell[     136] = 32'h0;  // 32'hf63bbeda;
    ram_cell[     137] = 32'h0;  // 32'h2e16b4d4;
    ram_cell[     138] = 32'h0;  // 32'h33693d73;
    ram_cell[     139] = 32'h0;  // 32'he7edc3bb;
    ram_cell[     140] = 32'h0;  // 32'h9cb6e286;
    ram_cell[     141] = 32'h0;  // 32'hd7205261;
    ram_cell[     142] = 32'h0;  // 32'h8e2cf6f5;
    ram_cell[     143] = 32'h0;  // 32'hfee8765a;
    ram_cell[     144] = 32'h0;  // 32'h00b07669;
    ram_cell[     145] = 32'h0;  // 32'h93488058;
    ram_cell[     146] = 32'h0;  // 32'hd42e7c44;
    ram_cell[     147] = 32'h0;  // 32'hc0a9a96d;
    ram_cell[     148] = 32'h0;  // 32'h1d5d9f6e;
    ram_cell[     149] = 32'h0;  // 32'hebf7e0d4;
    ram_cell[     150] = 32'h0;  // 32'h4c43aa0a;
    ram_cell[     151] = 32'h0;  // 32'h00680447;
    ram_cell[     152] = 32'h0;  // 32'h5c13b638;
    ram_cell[     153] = 32'h0;  // 32'h6ad5870c;
    ram_cell[     154] = 32'h0;  // 32'h854f64d7;
    ram_cell[     155] = 32'h0;  // 32'h95b3a5dd;
    ram_cell[     156] = 32'h0;  // 32'h0dc71199;
    ram_cell[     157] = 32'h0;  // 32'h3f8b45a1;
    ram_cell[     158] = 32'h0;  // 32'h1ec0ef0b;
    ram_cell[     159] = 32'h0;  // 32'hd5c99bf6;
    ram_cell[     160] = 32'h0;  // 32'hb7eb46fc;
    ram_cell[     161] = 32'h0;  // 32'h5ad07c52;
    ram_cell[     162] = 32'h0;  // 32'hfdaa9eca;
    ram_cell[     163] = 32'h0;  // 32'h0be8bb7b;
    ram_cell[     164] = 32'h0;  // 32'hf8cadf48;
    ram_cell[     165] = 32'h0;  // 32'h127e02b4;
    ram_cell[     166] = 32'h0;  // 32'h363edd9f;
    ram_cell[     167] = 32'h0;  // 32'ha9c0e82d;
    ram_cell[     168] = 32'h0;  // 32'h1334fea7;
    ram_cell[     169] = 32'h0;  // 32'hbcd13fd8;
    ram_cell[     170] = 32'h0;  // 32'h0f845869;
    ram_cell[     171] = 32'h0;  // 32'h6804b447;
    ram_cell[     172] = 32'h0;  // 32'h371c60e1;
    ram_cell[     173] = 32'h0;  // 32'h9b2e6349;
    ram_cell[     174] = 32'h0;  // 32'h57e4fb68;
    ram_cell[     175] = 32'h0;  // 32'h3f29fe33;
    ram_cell[     176] = 32'h0;  // 32'h1e9218a1;
    ram_cell[     177] = 32'h0;  // 32'hd8cf7574;
    ram_cell[     178] = 32'h0;  // 32'h3a54b80a;
    ram_cell[     179] = 32'h0;  // 32'h035dbe2b;
    ram_cell[     180] = 32'h0;  // 32'had565ea6;
    ram_cell[     181] = 32'h0;  // 32'h4b052072;
    ram_cell[     182] = 32'h0;  // 32'h179b5cf7;
    ram_cell[     183] = 32'h0;  // 32'h9af3abb6;
    ram_cell[     184] = 32'h0;  // 32'h86e46972;
    ram_cell[     185] = 32'h0;  // 32'h6d3bdee4;
    ram_cell[     186] = 32'h0;  // 32'hccddd93a;
    ram_cell[     187] = 32'h0;  // 32'hdf54d03b;
    ram_cell[     188] = 32'h0;  // 32'h28002bdc;
    ram_cell[     189] = 32'h0;  // 32'h4ddf9dec;
    ram_cell[     190] = 32'h0;  // 32'h0106b64f;
    ram_cell[     191] = 32'h0;  // 32'h62011113;
    ram_cell[     192] = 32'h0;  // 32'heac94584;
    ram_cell[     193] = 32'h0;  // 32'h28d375d2;
    ram_cell[     194] = 32'h0;  // 32'h46d82368;
    ram_cell[     195] = 32'h0;  // 32'hdabc7daf;
    ram_cell[     196] = 32'h0;  // 32'hfdad0898;
    ram_cell[     197] = 32'h0;  // 32'h709da868;
    ram_cell[     198] = 32'h0;  // 32'h7ca29683;
    ram_cell[     199] = 32'h0;  // 32'h167a2820;
    ram_cell[     200] = 32'h0;  // 32'hf6c6b6fc;
    ram_cell[     201] = 32'h0;  // 32'h277418fa;
    ram_cell[     202] = 32'h0;  // 32'h4e5f5eb5;
    ram_cell[     203] = 32'h0;  // 32'h8d274fd5;
    ram_cell[     204] = 32'h0;  // 32'h4080249e;
    ram_cell[     205] = 32'h0;  // 32'heeaa5cd9;
    ram_cell[     206] = 32'h0;  // 32'h0e99b45d;
    ram_cell[     207] = 32'h0;  // 32'h2fcecfee;
    ram_cell[     208] = 32'h0;  // 32'h42482da8;
    ram_cell[     209] = 32'h0;  // 32'h3a425038;
    ram_cell[     210] = 32'h0;  // 32'h48cd9664;
    ram_cell[     211] = 32'h0;  // 32'h32f5d3db;
    ram_cell[     212] = 32'h0;  // 32'hee312bd9;
    ram_cell[     213] = 32'h0;  // 32'h2bc940f1;
    ram_cell[     214] = 32'h0;  // 32'h37ee571d;
    ram_cell[     215] = 32'h0;  // 32'hb0b7981f;
    ram_cell[     216] = 32'h0;  // 32'hb445c73b;
    ram_cell[     217] = 32'h0;  // 32'h27d133d6;
    ram_cell[     218] = 32'h0;  // 32'hf74dd0fc;
    ram_cell[     219] = 32'h0;  // 32'h38edda28;
    ram_cell[     220] = 32'h0;  // 32'h262944f4;
    ram_cell[     221] = 32'h0;  // 32'hd06f078f;
    ram_cell[     222] = 32'h0;  // 32'h11cb35f7;
    ram_cell[     223] = 32'h0;  // 32'h6d0b475a;
    ram_cell[     224] = 32'h0;  // 32'h03ce3152;
    ram_cell[     225] = 32'h0;  // 32'h0fa0ad3b;
    ram_cell[     226] = 32'h0;  // 32'h5c28c288;
    ram_cell[     227] = 32'h0;  // 32'h3005b4de;
    ram_cell[     228] = 32'h0;  // 32'ha4cbd790;
    ram_cell[     229] = 32'h0;  // 32'hb367c55c;
    ram_cell[     230] = 32'h0;  // 32'hf74388f2;
    ram_cell[     231] = 32'h0;  // 32'ha1165ffa;
    ram_cell[     232] = 32'h0;  // 32'he56e64e3;
    ram_cell[     233] = 32'h0;  // 32'hee98e138;
    ram_cell[     234] = 32'h0;  // 32'ha79d183d;
    ram_cell[     235] = 32'h0;  // 32'h0dfa1f08;
    ram_cell[     236] = 32'h0;  // 32'h501b087d;
    ram_cell[     237] = 32'h0;  // 32'h73b7ef36;
    ram_cell[     238] = 32'h0;  // 32'h8e53ff63;
    ram_cell[     239] = 32'h0;  // 32'hd43e8280;
    ram_cell[     240] = 32'h0;  // 32'hefed07c1;
    ram_cell[     241] = 32'h0;  // 32'hcae8f612;
    ram_cell[     242] = 32'h0;  // 32'he6339baf;
    ram_cell[     243] = 32'h0;  // 32'h84f5b4a2;
    ram_cell[     244] = 32'h0;  // 32'h3d554028;
    ram_cell[     245] = 32'h0;  // 32'h49f12ac2;
    ram_cell[     246] = 32'h0;  // 32'h6e9a9d55;
    ram_cell[     247] = 32'h0;  // 32'hf4d90cc6;
    ram_cell[     248] = 32'h0;  // 32'h62978660;
    ram_cell[     249] = 32'h0;  // 32'h866eaab0;
    ram_cell[     250] = 32'h0;  // 32'h5a41f0da;
    ram_cell[     251] = 32'h0;  // 32'h1c3cf8c3;
    ram_cell[     252] = 32'h0;  // 32'h69e69661;
    ram_cell[     253] = 32'h0;  // 32'h03fc735a;
    ram_cell[     254] = 32'h0;  // 32'h890f17ef;
    ram_cell[     255] = 32'h0;  // 32'h96402147;
    // src matrix A
    ram_cell[     256] = 32'h79d54295;
    ram_cell[     257] = 32'h1be069a4;
    ram_cell[     258] = 32'h36a3234b;
    ram_cell[     259] = 32'h1a3e9280;
    ram_cell[     260] = 32'h71d06870;
    ram_cell[     261] = 32'hdeea0266;
    ram_cell[     262] = 32'h63aca52d;
    ram_cell[     263] = 32'h23a0d00d;
    ram_cell[     264] = 32'h33436186;
    ram_cell[     265] = 32'ha9b34353;
    ram_cell[     266] = 32'h12ba0d56;
    ram_cell[     267] = 32'h5b40d795;
    ram_cell[     268] = 32'hf1a05c49;
    ram_cell[     269] = 32'hedafd7ac;
    ram_cell[     270] = 32'hefef2311;
    ram_cell[     271] = 32'hee0b2090;
    ram_cell[     272] = 32'h10cf1a6d;
    ram_cell[     273] = 32'hd31a8c9e;
    ram_cell[     274] = 32'h27fc9fd0;
    ram_cell[     275] = 32'h87a5cd61;
    ram_cell[     276] = 32'ha4058cdc;
    ram_cell[     277] = 32'hd0840424;
    ram_cell[     278] = 32'h6ea77c50;
    ram_cell[     279] = 32'hb8bcaff8;
    ram_cell[     280] = 32'h3ddd7cfd;
    ram_cell[     281] = 32'h4a023bbe;
    ram_cell[     282] = 32'h0d5d282b;
    ram_cell[     283] = 32'hbfb99f55;
    ram_cell[     284] = 32'h2b95b8b3;
    ram_cell[     285] = 32'h3adf9ed1;
    ram_cell[     286] = 32'h1cdef4a8;
    ram_cell[     287] = 32'hd8e684c2;
    ram_cell[     288] = 32'h1243dced;
    ram_cell[     289] = 32'h12731193;
    ram_cell[     290] = 32'hb4e83b95;
    ram_cell[     291] = 32'h62b21b3c;
    ram_cell[     292] = 32'h34be39ec;
    ram_cell[     293] = 32'hc89cf3d8;
    ram_cell[     294] = 32'hebe8f2bd;
    ram_cell[     295] = 32'h8e98606f;
    ram_cell[     296] = 32'h871cb9c0;
    ram_cell[     297] = 32'h4964c036;
    ram_cell[     298] = 32'h07e2e776;
    ram_cell[     299] = 32'h392e0988;
    ram_cell[     300] = 32'h82b2ec63;
    ram_cell[     301] = 32'h23e0458b;
    ram_cell[     302] = 32'h20b370d8;
    ram_cell[     303] = 32'h23e20ca3;
    ram_cell[     304] = 32'hddb57cbd;
    ram_cell[     305] = 32'h2d827630;
    ram_cell[     306] = 32'h884f43a7;
    ram_cell[     307] = 32'hfe17a387;
    ram_cell[     308] = 32'h03009367;
    ram_cell[     309] = 32'h49743d9d;
    ram_cell[     310] = 32'h639db8f2;
    ram_cell[     311] = 32'he16dcd80;
    ram_cell[     312] = 32'h97d43917;
    ram_cell[     313] = 32'h287bceb1;
    ram_cell[     314] = 32'h42de7e5b;
    ram_cell[     315] = 32'hfb7ac563;
    ram_cell[     316] = 32'h55be7ed3;
    ram_cell[     317] = 32'hd4af0cdb;
    ram_cell[     318] = 32'h3d0d2146;
    ram_cell[     319] = 32'ha86e2a08;
    ram_cell[     320] = 32'h80f40b8f;
    ram_cell[     321] = 32'h018f7d4f;
    ram_cell[     322] = 32'h17c7fe62;
    ram_cell[     323] = 32'hf6f8ccfe;
    ram_cell[     324] = 32'h099ae7d3;
    ram_cell[     325] = 32'h522b4fea;
    ram_cell[     326] = 32'ha99cf3c6;
    ram_cell[     327] = 32'hab931318;
    ram_cell[     328] = 32'h4d5df9b0;
    ram_cell[     329] = 32'ha1e7c335;
    ram_cell[     330] = 32'h4f4beba8;
    ram_cell[     331] = 32'h7c8cc509;
    ram_cell[     332] = 32'hd5cf1a8c;
    ram_cell[     333] = 32'hc7560e49;
    ram_cell[     334] = 32'h4b01690b;
    ram_cell[     335] = 32'h3732382f;
    ram_cell[     336] = 32'hb2496e2e;
    ram_cell[     337] = 32'hcc46f159;
    ram_cell[     338] = 32'h6870e534;
    ram_cell[     339] = 32'he448b3ae;
    ram_cell[     340] = 32'hf248281a;
    ram_cell[     341] = 32'hd94f8e7a;
    ram_cell[     342] = 32'hf4bb2a3a;
    ram_cell[     343] = 32'h27da72ad;
    ram_cell[     344] = 32'h46bab040;
    ram_cell[     345] = 32'h2347c41f;
    ram_cell[     346] = 32'h912e5e9e;
    ram_cell[     347] = 32'hd9c04049;
    ram_cell[     348] = 32'h39071954;
    ram_cell[     349] = 32'h744c788c;
    ram_cell[     350] = 32'h3144abb3;
    ram_cell[     351] = 32'h2efb405c;
    ram_cell[     352] = 32'hee60adca;
    ram_cell[     353] = 32'h09e95a1a;
    ram_cell[     354] = 32'h85609cf7;
    ram_cell[     355] = 32'hea4a9be0;
    ram_cell[     356] = 32'h8c1b41b3;
    ram_cell[     357] = 32'h1ccefa13;
    ram_cell[     358] = 32'h793e0df1;
    ram_cell[     359] = 32'h09a70ee4;
    ram_cell[     360] = 32'h4ba37600;
    ram_cell[     361] = 32'hf2bd3d5c;
    ram_cell[     362] = 32'h36eaef8f;
    ram_cell[     363] = 32'h1ee94ffb;
    ram_cell[     364] = 32'h785b3af9;
    ram_cell[     365] = 32'hfb883206;
    ram_cell[     366] = 32'h84e73a18;
    ram_cell[     367] = 32'hd0c0c056;
    ram_cell[     368] = 32'hf3da9979;
    ram_cell[     369] = 32'hb2ce883d;
    ram_cell[     370] = 32'h7644bc9d;
    ram_cell[     371] = 32'h3311c2dd;
    ram_cell[     372] = 32'h5c5302b8;
    ram_cell[     373] = 32'h11e52731;
    ram_cell[     374] = 32'he796c57e;
    ram_cell[     375] = 32'h95da0c42;
    ram_cell[     376] = 32'hda6388da;
    ram_cell[     377] = 32'he7accc2a;
    ram_cell[     378] = 32'ha918527d;
    ram_cell[     379] = 32'hf8fad089;
    ram_cell[     380] = 32'hf1c1b064;
    ram_cell[     381] = 32'hc27be517;
    ram_cell[     382] = 32'h73632b3d;
    ram_cell[     383] = 32'h2df4b972;
    ram_cell[     384] = 32'h786ee65b;
    ram_cell[     385] = 32'ha210f5d6;
    ram_cell[     386] = 32'he18020af;
    ram_cell[     387] = 32'h04c56e9d;
    ram_cell[     388] = 32'hbcd31e5c;
    ram_cell[     389] = 32'hd08d1023;
    ram_cell[     390] = 32'ha874b755;
    ram_cell[     391] = 32'hcc92d227;
    ram_cell[     392] = 32'h984e1a4e;
    ram_cell[     393] = 32'hd45a1c3d;
    ram_cell[     394] = 32'h6ba88c2b;
    ram_cell[     395] = 32'h48b3372b;
    ram_cell[     396] = 32'h408db575;
    ram_cell[     397] = 32'h8bf1bd98;
    ram_cell[     398] = 32'h77708fa1;
    ram_cell[     399] = 32'h7ab3da20;
    ram_cell[     400] = 32'hb573e2dd;
    ram_cell[     401] = 32'h037fd4aa;
    ram_cell[     402] = 32'h1c88e07c;
    ram_cell[     403] = 32'h79374a81;
    ram_cell[     404] = 32'h46d1b1c0;
    ram_cell[     405] = 32'h05e851f1;
    ram_cell[     406] = 32'hc3f19b19;
    ram_cell[     407] = 32'h72f98da0;
    ram_cell[     408] = 32'h36495b67;
    ram_cell[     409] = 32'h14ae8355;
    ram_cell[     410] = 32'h9554ad24;
    ram_cell[     411] = 32'h150ff773;
    ram_cell[     412] = 32'h6a2aec6b;
    ram_cell[     413] = 32'h78e653d8;
    ram_cell[     414] = 32'h4d4d9e9e;
    ram_cell[     415] = 32'h14970da1;
    ram_cell[     416] = 32'h63c40616;
    ram_cell[     417] = 32'hb727856a;
    ram_cell[     418] = 32'h7b41c6b1;
    ram_cell[     419] = 32'h66cae935;
    ram_cell[     420] = 32'h9220afe1;
    ram_cell[     421] = 32'hbf935a70;
    ram_cell[     422] = 32'hd94214ce;
    ram_cell[     423] = 32'hc95f7e46;
    ram_cell[     424] = 32'hd3003fd4;
    ram_cell[     425] = 32'h2c915eb1;
    ram_cell[     426] = 32'hf5bcaac5;
    ram_cell[     427] = 32'hfafc9742;
    ram_cell[     428] = 32'hbde0775c;
    ram_cell[     429] = 32'h8c9185a3;
    ram_cell[     430] = 32'ha44a1115;
    ram_cell[     431] = 32'hc1f3ad2e;
    ram_cell[     432] = 32'hb0754d0d;
    ram_cell[     433] = 32'hcf79b966;
    ram_cell[     434] = 32'h33883d4a;
    ram_cell[     435] = 32'h6b4a4d31;
    ram_cell[     436] = 32'h230f4533;
    ram_cell[     437] = 32'h1c383b3a;
    ram_cell[     438] = 32'hf7513af1;
    ram_cell[     439] = 32'hefd4711d;
    ram_cell[     440] = 32'h061d6e83;
    ram_cell[     441] = 32'h03b496f7;
    ram_cell[     442] = 32'hb6630e7f;
    ram_cell[     443] = 32'hb772a29f;
    ram_cell[     444] = 32'h750efbcd;
    ram_cell[     445] = 32'hccc622f7;
    ram_cell[     446] = 32'h00f3aebe;
    ram_cell[     447] = 32'h7c7da21d;
    ram_cell[     448] = 32'h03814991;
    ram_cell[     449] = 32'h45146f22;
    ram_cell[     450] = 32'h59e2cb81;
    ram_cell[     451] = 32'hd98b0f7d;
    ram_cell[     452] = 32'h8c96b03b;
    ram_cell[     453] = 32'he646f709;
    ram_cell[     454] = 32'h038c8634;
    ram_cell[     455] = 32'h22161718;
    ram_cell[     456] = 32'hb0aca2f2;
    ram_cell[     457] = 32'h8b2e5175;
    ram_cell[     458] = 32'h23282405;
    ram_cell[     459] = 32'h2c676ee4;
    ram_cell[     460] = 32'hb301c550;
    ram_cell[     461] = 32'h5164f135;
    ram_cell[     462] = 32'h575d5886;
    ram_cell[     463] = 32'hff852cda;
    ram_cell[     464] = 32'h2faa3c9e;
    ram_cell[     465] = 32'h7d116252;
    ram_cell[     466] = 32'ha1c4d920;
    ram_cell[     467] = 32'h463b7b29;
    ram_cell[     468] = 32'hd9dde829;
    ram_cell[     469] = 32'h12c02bd9;
    ram_cell[     470] = 32'hf87a4113;
    ram_cell[     471] = 32'h7439eea3;
    ram_cell[     472] = 32'h933e3a71;
    ram_cell[     473] = 32'hbe00b8db;
    ram_cell[     474] = 32'hadfeeebf;
    ram_cell[     475] = 32'hc5f81c39;
    ram_cell[     476] = 32'h0d97461c;
    ram_cell[     477] = 32'h7d296e69;
    ram_cell[     478] = 32'h7068dc82;
    ram_cell[     479] = 32'hc99811e7;
    ram_cell[     480] = 32'h2c241e36;
    ram_cell[     481] = 32'hef405331;
    ram_cell[     482] = 32'h91c10cc6;
    ram_cell[     483] = 32'hc4b36740;
    ram_cell[     484] = 32'hb517f873;
    ram_cell[     485] = 32'h14848b27;
    ram_cell[     486] = 32'hf076f077;
    ram_cell[     487] = 32'h938a39fc;
    ram_cell[     488] = 32'h3f98b4f9;
    ram_cell[     489] = 32'h798d1caf;
    ram_cell[     490] = 32'h243e64bc;
    ram_cell[     491] = 32'h2959684c;
    ram_cell[     492] = 32'hd59f8fec;
    ram_cell[     493] = 32'hdb246ae8;
    ram_cell[     494] = 32'h97986028;
    ram_cell[     495] = 32'hf71f596e;
    ram_cell[     496] = 32'h34b62781;
    ram_cell[     497] = 32'h5f3444c2;
    ram_cell[     498] = 32'ha9e4842c;
    ram_cell[     499] = 32'h74650ea8;
    ram_cell[     500] = 32'h537f67e9;
    ram_cell[     501] = 32'h79e228b7;
    ram_cell[     502] = 32'hc4fdf28d;
    ram_cell[     503] = 32'hb768bf50;
    ram_cell[     504] = 32'h31311d52;
    ram_cell[     505] = 32'h2800e732;
    ram_cell[     506] = 32'hc1138dbb;
    ram_cell[     507] = 32'h560e9408;
    ram_cell[     508] = 32'heeebecef;
    ram_cell[     509] = 32'h8d1d3315;
    ram_cell[     510] = 32'hcd1d02aa;
    ram_cell[     511] = 32'hedad6e3f;
    // src matrix B
    ram_cell[     512] = 32'h8a0195c4;
    ram_cell[     513] = 32'h5fb9e47d;
    ram_cell[     514] = 32'h8f5d40fa;
    ram_cell[     515] = 32'h79f89965;
    ram_cell[     516] = 32'h4686ca68;
    ram_cell[     517] = 32'h96941d8c;
    ram_cell[     518] = 32'h7aa351cc;
    ram_cell[     519] = 32'h211d3ae7;
    ram_cell[     520] = 32'he202d327;
    ram_cell[     521] = 32'h41ccae66;
    ram_cell[     522] = 32'h4650c660;
    ram_cell[     523] = 32'ha878d8a2;
    ram_cell[     524] = 32'h44ee38ea;
    ram_cell[     525] = 32'h08cd832e;
    ram_cell[     526] = 32'hef9b78ee;
    ram_cell[     527] = 32'h00fdb56e;
    ram_cell[     528] = 32'haf3e2401;
    ram_cell[     529] = 32'h8b2652db;
    ram_cell[     530] = 32'h51a7dc7a;
    ram_cell[     531] = 32'h2a7ca794;
    ram_cell[     532] = 32'hc28928f6;
    ram_cell[     533] = 32'h0ef8c9ec;
    ram_cell[     534] = 32'h5c8e4407;
    ram_cell[     535] = 32'h4a5ae8fe;
    ram_cell[     536] = 32'h21e6dc85;
    ram_cell[     537] = 32'h92b9dffd;
    ram_cell[     538] = 32'hfe18aa0c;
    ram_cell[     539] = 32'hb252435a;
    ram_cell[     540] = 32'h89c18377;
    ram_cell[     541] = 32'h145980fe;
    ram_cell[     542] = 32'h2de64f9f;
    ram_cell[     543] = 32'h32c48c0d;
    ram_cell[     544] = 32'h2b3ab5fb;
    ram_cell[     545] = 32'h9db9ee37;
    ram_cell[     546] = 32'h2ef63a03;
    ram_cell[     547] = 32'hd7caa125;
    ram_cell[     548] = 32'heca5f9d4;
    ram_cell[     549] = 32'h5c16a915;
    ram_cell[     550] = 32'hf250bac1;
    ram_cell[     551] = 32'hf09b3ea1;
    ram_cell[     552] = 32'hbd60ef7d;
    ram_cell[     553] = 32'h27d786ba;
    ram_cell[     554] = 32'h17318d27;
    ram_cell[     555] = 32'hc7d3a447;
    ram_cell[     556] = 32'h5433a304;
    ram_cell[     557] = 32'h186e238d;
    ram_cell[     558] = 32'h4efde05a;
    ram_cell[     559] = 32'h148cc8c9;
    ram_cell[     560] = 32'hec040f1b;
    ram_cell[     561] = 32'h415fc0c4;
    ram_cell[     562] = 32'h10696454;
    ram_cell[     563] = 32'h7175ee11;
    ram_cell[     564] = 32'ha3208324;
    ram_cell[     565] = 32'h4a9643ba;
    ram_cell[     566] = 32'hd129f69a;
    ram_cell[     567] = 32'h14568e30;
    ram_cell[     568] = 32'haf0bb47c;
    ram_cell[     569] = 32'h4adc93d1;
    ram_cell[     570] = 32'hb4f67fe2;
    ram_cell[     571] = 32'h690268ee;
    ram_cell[     572] = 32'h6f9dc12b;
    ram_cell[     573] = 32'h85ac13cc;
    ram_cell[     574] = 32'h9e86e18f;
    ram_cell[     575] = 32'hf2794986;
    ram_cell[     576] = 32'h36292b20;
    ram_cell[     577] = 32'hf9b10a0d;
    ram_cell[     578] = 32'h912e60da;
    ram_cell[     579] = 32'h163fb4c4;
    ram_cell[     580] = 32'h90c0f067;
    ram_cell[     581] = 32'haa38483c;
    ram_cell[     582] = 32'h68a13ce2;
    ram_cell[     583] = 32'h41370345;
    ram_cell[     584] = 32'h10ca1b25;
    ram_cell[     585] = 32'h4a9f9224;
    ram_cell[     586] = 32'h1f8f8ab4;
    ram_cell[     587] = 32'h03432712;
    ram_cell[     588] = 32'he1ded2b6;
    ram_cell[     589] = 32'h071037c2;
    ram_cell[     590] = 32'hb60686b0;
    ram_cell[     591] = 32'h032adabc;
    ram_cell[     592] = 32'h6838b6b5;
    ram_cell[     593] = 32'he11c514e;
    ram_cell[     594] = 32'h0e0a0ffb;
    ram_cell[     595] = 32'he550a51e;
    ram_cell[     596] = 32'h48c03574;
    ram_cell[     597] = 32'h88535cf1;
    ram_cell[     598] = 32'hd377cfe0;
    ram_cell[     599] = 32'he235c4aa;
    ram_cell[     600] = 32'h3c04ecbe;
    ram_cell[     601] = 32'hf6497303;
    ram_cell[     602] = 32'h57cad88f;
    ram_cell[     603] = 32'h0c691f21;
    ram_cell[     604] = 32'hbc87150c;
    ram_cell[     605] = 32'h8dba9cb5;
    ram_cell[     606] = 32'h0d6ba409;
    ram_cell[     607] = 32'h7dbc97e1;
    ram_cell[     608] = 32'h1ea80e41;
    ram_cell[     609] = 32'h32fdf600;
    ram_cell[     610] = 32'h930a9342;
    ram_cell[     611] = 32'h5981ce98;
    ram_cell[     612] = 32'h1fc9f336;
    ram_cell[     613] = 32'h0aaec863;
    ram_cell[     614] = 32'hdeaf8bdc;
    ram_cell[     615] = 32'hb442153b;
    ram_cell[     616] = 32'h74213e2b;
    ram_cell[     617] = 32'h885f193e;
    ram_cell[     618] = 32'hfe346157;
    ram_cell[     619] = 32'h430980e4;
    ram_cell[     620] = 32'h07344026;
    ram_cell[     621] = 32'h83abbb5a;
    ram_cell[     622] = 32'h979584b1;
    ram_cell[     623] = 32'h0c899ef8;
    ram_cell[     624] = 32'h64addefe;
    ram_cell[     625] = 32'hfcfb96b2;
    ram_cell[     626] = 32'h3f54f04a;
    ram_cell[     627] = 32'h4683ed81;
    ram_cell[     628] = 32'hd2bfea22;
    ram_cell[     629] = 32'hbc3ee099;
    ram_cell[     630] = 32'h01e3152e;
    ram_cell[     631] = 32'h024ca82b;
    ram_cell[     632] = 32'h12bf3541;
    ram_cell[     633] = 32'heafea7ea;
    ram_cell[     634] = 32'h1ecc405b;
    ram_cell[     635] = 32'hd4473e4e;
    ram_cell[     636] = 32'h120e99f4;
    ram_cell[     637] = 32'h4d1733a4;
    ram_cell[     638] = 32'h3d19da30;
    ram_cell[     639] = 32'h412861a3;
    ram_cell[     640] = 32'h421f90b1;
    ram_cell[     641] = 32'h430165cf;
    ram_cell[     642] = 32'h3d208f00;
    ram_cell[     643] = 32'h68c75ecb;
    ram_cell[     644] = 32'hc3264363;
    ram_cell[     645] = 32'hfdd4047a;
    ram_cell[     646] = 32'hc60c520e;
    ram_cell[     647] = 32'h4d675b30;
    ram_cell[     648] = 32'hcc025c35;
    ram_cell[     649] = 32'h084b0287;
    ram_cell[     650] = 32'h39310515;
    ram_cell[     651] = 32'hca75fcb7;
    ram_cell[     652] = 32'hc7b655c6;
    ram_cell[     653] = 32'h396f3d1e;
    ram_cell[     654] = 32'h28a5075e;
    ram_cell[     655] = 32'h1277cc77;
    ram_cell[     656] = 32'h168723a0;
    ram_cell[     657] = 32'h6d02461e;
    ram_cell[     658] = 32'h1628d3d5;
    ram_cell[     659] = 32'hf46b1391;
    ram_cell[     660] = 32'h031ddc44;
    ram_cell[     661] = 32'hf8342e26;
    ram_cell[     662] = 32'h0d84a129;
    ram_cell[     663] = 32'h18974a76;
    ram_cell[     664] = 32'hfd9938b5;
    ram_cell[     665] = 32'ha440620d;
    ram_cell[     666] = 32'h1c69e3d0;
    ram_cell[     667] = 32'hee4c7af4;
    ram_cell[     668] = 32'hed71f1cc;
    ram_cell[     669] = 32'hc0795245;
    ram_cell[     670] = 32'hf4c2e6f4;
    ram_cell[     671] = 32'h27f674eb;
    ram_cell[     672] = 32'h0751f9fd;
    ram_cell[     673] = 32'h64597bad;
    ram_cell[     674] = 32'ha5cd41f0;
    ram_cell[     675] = 32'h6e2ba1ec;
    ram_cell[     676] = 32'hf36918c6;
    ram_cell[     677] = 32'hb6d4e5bf;
    ram_cell[     678] = 32'he830bc9c;
    ram_cell[     679] = 32'hcad2b58f;
    ram_cell[     680] = 32'h9ae217c0;
    ram_cell[     681] = 32'h0f49841b;
    ram_cell[     682] = 32'hf10913a4;
    ram_cell[     683] = 32'h3c62f072;
    ram_cell[     684] = 32'hd5f58e8a;
    ram_cell[     685] = 32'hc54595cb;
    ram_cell[     686] = 32'h0b891c41;
    ram_cell[     687] = 32'he4794962;
    ram_cell[     688] = 32'h7ef76217;
    ram_cell[     689] = 32'h21155611;
    ram_cell[     690] = 32'hc35bc223;
    ram_cell[     691] = 32'h7698c169;
    ram_cell[     692] = 32'h9c8eae93;
    ram_cell[     693] = 32'h9db3835a;
    ram_cell[     694] = 32'haaac9193;
    ram_cell[     695] = 32'h24a3e0d9;
    ram_cell[     696] = 32'h3174cd1d;
    ram_cell[     697] = 32'he016ac96;
    ram_cell[     698] = 32'h917c166b;
    ram_cell[     699] = 32'h5c50e46c;
    ram_cell[     700] = 32'hdf6b9628;
    ram_cell[     701] = 32'h26a73ba4;
    ram_cell[     702] = 32'h4cd010f4;
    ram_cell[     703] = 32'h8c975d06;
    ram_cell[     704] = 32'hbf54cbc2;
    ram_cell[     705] = 32'h9572be75;
    ram_cell[     706] = 32'h4812222d;
    ram_cell[     707] = 32'h7ad1e9cf;
    ram_cell[     708] = 32'h5d4eea37;
    ram_cell[     709] = 32'hcd2c0aee;
    ram_cell[     710] = 32'he7af049e;
    ram_cell[     711] = 32'h84a32b98;
    ram_cell[     712] = 32'hdec005d2;
    ram_cell[     713] = 32'h2a5f55d7;
    ram_cell[     714] = 32'h4f62c4a3;
    ram_cell[     715] = 32'h401782ce;
    ram_cell[     716] = 32'h577b4d00;
    ram_cell[     717] = 32'h57ab1a86;
    ram_cell[     718] = 32'hafbef499;
    ram_cell[     719] = 32'h8b24d306;
    ram_cell[     720] = 32'h09c48018;
    ram_cell[     721] = 32'h5a04e1e8;
    ram_cell[     722] = 32'h11227771;
    ram_cell[     723] = 32'hefe56c75;
    ram_cell[     724] = 32'hcb90c879;
    ram_cell[     725] = 32'hc38197ef;
    ram_cell[     726] = 32'h70a9bf55;
    ram_cell[     727] = 32'h9e3da936;
    ram_cell[     728] = 32'h846db0f4;
    ram_cell[     729] = 32'he7c83434;
    ram_cell[     730] = 32'h2b45acd9;
    ram_cell[     731] = 32'h7aaf3297;
    ram_cell[     732] = 32'h2ac618ff;
    ram_cell[     733] = 32'h42b6f211;
    ram_cell[     734] = 32'h2b3c898e;
    ram_cell[     735] = 32'h072867df;
    ram_cell[     736] = 32'h6361f849;
    ram_cell[     737] = 32'hb0d70f45;
    ram_cell[     738] = 32'hc1ad6d61;
    ram_cell[     739] = 32'h54e96887;
    ram_cell[     740] = 32'hc7eae2f6;
    ram_cell[     741] = 32'hd1cab1ad;
    ram_cell[     742] = 32'hfaa813ac;
    ram_cell[     743] = 32'h66f362be;
    ram_cell[     744] = 32'h95cab2a0;
    ram_cell[     745] = 32'hdc66ecbd;
    ram_cell[     746] = 32'hb05c7c03;
    ram_cell[     747] = 32'h3047c419;
    ram_cell[     748] = 32'h8d3f0e89;
    ram_cell[     749] = 32'h897e6f39;
    ram_cell[     750] = 32'h2ac2140e;
    ram_cell[     751] = 32'h7a91823c;
    ram_cell[     752] = 32'h630c9228;
    ram_cell[     753] = 32'h04474a2a;
    ram_cell[     754] = 32'h99510294;
    ram_cell[     755] = 32'h9c0f4277;
    ram_cell[     756] = 32'hdf86e28b;
    ram_cell[     757] = 32'h24c26c5a;
    ram_cell[     758] = 32'h317815fa;
    ram_cell[     759] = 32'h8c092f7c;
    ram_cell[     760] = 32'h57f236ed;
    ram_cell[     761] = 32'h702c00b9;
    ram_cell[     762] = 32'ha18d9b1c;
    ram_cell[     763] = 32'h640588c9;
    ram_cell[     764] = 32'h4c26658a;
    ram_cell[     765] = 32'h9ac0b7eb;
    ram_cell[     766] = 32'h22921491;
    ram_cell[     767] = 32'hd4e69615;
end

endmodule

