
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h1a6333ec;
    ram_cell[       1] = 32'h0;  // 32'hf38d8cf6;
    ram_cell[       2] = 32'h0;  // 32'h9bd3c175;
    ram_cell[       3] = 32'h0;  // 32'h45eafa1a;
    ram_cell[       4] = 32'h0;  // 32'h8a850bdc;
    ram_cell[       5] = 32'h0;  // 32'hba58a66b;
    ram_cell[       6] = 32'h0;  // 32'hf684c846;
    ram_cell[       7] = 32'h0;  // 32'h61a736c1;
    ram_cell[       8] = 32'h0;  // 32'h42b3f444;
    ram_cell[       9] = 32'h0;  // 32'h44dbcf10;
    ram_cell[      10] = 32'h0;  // 32'hff2ce9c0;
    ram_cell[      11] = 32'h0;  // 32'h93d70847;
    ram_cell[      12] = 32'h0;  // 32'h90d9230b;
    ram_cell[      13] = 32'h0;  // 32'hb4536433;
    ram_cell[      14] = 32'h0;  // 32'h376082b8;
    ram_cell[      15] = 32'h0;  // 32'h4ed62c79;
    ram_cell[      16] = 32'h0;  // 32'h2204adc9;
    ram_cell[      17] = 32'h0;  // 32'h8e29d740;
    ram_cell[      18] = 32'h0;  // 32'h7f33cd64;
    ram_cell[      19] = 32'h0;  // 32'ha335621f;
    ram_cell[      20] = 32'h0;  // 32'h72c44bb3;
    ram_cell[      21] = 32'h0;  // 32'h600a0008;
    ram_cell[      22] = 32'h0;  // 32'h97b5e2ca;
    ram_cell[      23] = 32'h0;  // 32'h2243f443;
    ram_cell[      24] = 32'h0;  // 32'h58c1151e;
    ram_cell[      25] = 32'h0;  // 32'hc18f07b2;
    ram_cell[      26] = 32'h0;  // 32'h7fe3f20e;
    ram_cell[      27] = 32'h0;  // 32'hf5b76114;
    ram_cell[      28] = 32'h0;  // 32'ha58831fe;
    ram_cell[      29] = 32'h0;  // 32'h5200e37d;
    ram_cell[      30] = 32'h0;  // 32'hd9215b54;
    ram_cell[      31] = 32'h0;  // 32'h7f8f6b33;
    ram_cell[      32] = 32'h0;  // 32'h5284dd13;
    ram_cell[      33] = 32'h0;  // 32'hefeb9e66;
    ram_cell[      34] = 32'h0;  // 32'hce20e173;
    ram_cell[      35] = 32'h0;  // 32'hda03a825;
    ram_cell[      36] = 32'h0;  // 32'h98bb372d;
    ram_cell[      37] = 32'h0;  // 32'hee6f5e15;
    ram_cell[      38] = 32'h0;  // 32'hfc66a3da;
    ram_cell[      39] = 32'h0;  // 32'h9626b940;
    ram_cell[      40] = 32'h0;  // 32'hd70a5bb8;
    ram_cell[      41] = 32'h0;  // 32'h03e7aed4;
    ram_cell[      42] = 32'h0;  // 32'h6711fc6a;
    ram_cell[      43] = 32'h0;  // 32'hd546ae2d;
    ram_cell[      44] = 32'h0;  // 32'hf809534d;
    ram_cell[      45] = 32'h0;  // 32'h2737de14;
    ram_cell[      46] = 32'h0;  // 32'h05950431;
    ram_cell[      47] = 32'h0;  // 32'hccf70a2b;
    ram_cell[      48] = 32'h0;  // 32'h5f10e577;
    ram_cell[      49] = 32'h0;  // 32'h04486e49;
    ram_cell[      50] = 32'h0;  // 32'h61a10ec4;
    ram_cell[      51] = 32'h0;  // 32'h914b8f7e;
    ram_cell[      52] = 32'h0;  // 32'h53d76b9c;
    ram_cell[      53] = 32'h0;  // 32'h97377327;
    ram_cell[      54] = 32'h0;  // 32'h55e91095;
    ram_cell[      55] = 32'h0;  // 32'ha3c6f0fe;
    ram_cell[      56] = 32'h0;  // 32'h2968c9f6;
    ram_cell[      57] = 32'h0;  // 32'h68a52a7b;
    ram_cell[      58] = 32'h0;  // 32'h112cf5a7;
    ram_cell[      59] = 32'h0;  // 32'heae51c43;
    ram_cell[      60] = 32'h0;  // 32'hc137e68d;
    ram_cell[      61] = 32'h0;  // 32'h68c463cd;
    ram_cell[      62] = 32'h0;  // 32'hb964d2c5;
    ram_cell[      63] = 32'h0;  // 32'hcdf715f3;
    ram_cell[      64] = 32'h0;  // 32'hd8a75424;
    ram_cell[      65] = 32'h0;  // 32'hfbbd116c;
    ram_cell[      66] = 32'h0;  // 32'hfa5bcb1d;
    ram_cell[      67] = 32'h0;  // 32'h80eae2e9;
    ram_cell[      68] = 32'h0;  // 32'h8fbf141c;
    ram_cell[      69] = 32'h0;  // 32'h0e7d0a50;
    ram_cell[      70] = 32'h0;  // 32'hcb07af77;
    ram_cell[      71] = 32'h0;  // 32'h0252437a;
    ram_cell[      72] = 32'h0;  // 32'h6640cb7b;
    ram_cell[      73] = 32'h0;  // 32'hd39a30ae;
    ram_cell[      74] = 32'h0;  // 32'hc99ca3f5;
    ram_cell[      75] = 32'h0;  // 32'h40a48817;
    ram_cell[      76] = 32'h0;  // 32'h7c5d91dc;
    ram_cell[      77] = 32'h0;  // 32'hc076e3dc;
    ram_cell[      78] = 32'h0;  // 32'h20fa098e;
    ram_cell[      79] = 32'h0;  // 32'hab472fdf;
    ram_cell[      80] = 32'h0;  // 32'h844df0c7;
    ram_cell[      81] = 32'h0;  // 32'h106fceb2;
    ram_cell[      82] = 32'h0;  // 32'h1d098394;
    ram_cell[      83] = 32'h0;  // 32'hbc9acb00;
    ram_cell[      84] = 32'h0;  // 32'h6489af03;
    ram_cell[      85] = 32'h0;  // 32'hdfd47c41;
    ram_cell[      86] = 32'h0;  // 32'hc468e349;
    ram_cell[      87] = 32'h0;  // 32'h529d1bab;
    ram_cell[      88] = 32'h0;  // 32'h205a907f;
    ram_cell[      89] = 32'h0;  // 32'h42af54ec;
    ram_cell[      90] = 32'h0;  // 32'h0e887d7e;
    ram_cell[      91] = 32'h0;  // 32'hd9e00bc6;
    ram_cell[      92] = 32'h0;  // 32'hbe4fb9ad;
    ram_cell[      93] = 32'h0;  // 32'h55ac2c2c;
    ram_cell[      94] = 32'h0;  // 32'he8f16059;
    ram_cell[      95] = 32'h0;  // 32'h807f6f04;
    ram_cell[      96] = 32'h0;  // 32'h7f437102;
    ram_cell[      97] = 32'h0;  // 32'h632d20f9;
    ram_cell[      98] = 32'h0;  // 32'hb8d37dbb;
    ram_cell[      99] = 32'h0;  // 32'h640e434c;
    ram_cell[     100] = 32'h0;  // 32'h3d46f03d;
    ram_cell[     101] = 32'h0;  // 32'he23f936a;
    ram_cell[     102] = 32'h0;  // 32'h3dec3234;
    ram_cell[     103] = 32'h0;  // 32'h2b6948b9;
    ram_cell[     104] = 32'h0;  // 32'h75ef0a0a;
    ram_cell[     105] = 32'h0;  // 32'hb41ec709;
    ram_cell[     106] = 32'h0;  // 32'hd20bb4f8;
    ram_cell[     107] = 32'h0;  // 32'h6f27de4b;
    ram_cell[     108] = 32'h0;  // 32'h4f147007;
    ram_cell[     109] = 32'h0;  // 32'hd6806702;
    ram_cell[     110] = 32'h0;  // 32'hd7a62791;
    ram_cell[     111] = 32'h0;  // 32'h9e8aa4e4;
    ram_cell[     112] = 32'h0;  // 32'hfbfdadbf;
    ram_cell[     113] = 32'h0;  // 32'hecc9e2de;
    ram_cell[     114] = 32'h0;  // 32'hd1dd9129;
    ram_cell[     115] = 32'h0;  // 32'hf38393af;
    ram_cell[     116] = 32'h0;  // 32'h766ae928;
    ram_cell[     117] = 32'h0;  // 32'hc5db1128;
    ram_cell[     118] = 32'h0;  // 32'hb50ab20f;
    ram_cell[     119] = 32'h0;  // 32'hf6287778;
    ram_cell[     120] = 32'h0;  // 32'ha4a3609c;
    ram_cell[     121] = 32'h0;  // 32'h8ac40568;
    ram_cell[     122] = 32'h0;  // 32'ha8baa8b6;
    ram_cell[     123] = 32'h0;  // 32'hf0909b46;
    ram_cell[     124] = 32'h0;  // 32'h4b7c34ea;
    ram_cell[     125] = 32'h0;  // 32'hae07d6a1;
    ram_cell[     126] = 32'h0;  // 32'h6cf0aab6;
    ram_cell[     127] = 32'h0;  // 32'hb8ae2a94;
    ram_cell[     128] = 32'h0;  // 32'h75caf870;
    ram_cell[     129] = 32'h0;  // 32'h59f98694;
    ram_cell[     130] = 32'h0;  // 32'h16562ddc;
    ram_cell[     131] = 32'h0;  // 32'he5e6f4b4;
    ram_cell[     132] = 32'h0;  // 32'h5f00179f;
    ram_cell[     133] = 32'h0;  // 32'h8cc0bcf3;
    ram_cell[     134] = 32'h0;  // 32'h5bf8c243;
    ram_cell[     135] = 32'h0;  // 32'h431430bf;
    ram_cell[     136] = 32'h0;  // 32'h5df72a9e;
    ram_cell[     137] = 32'h0;  // 32'hf3a4e611;
    ram_cell[     138] = 32'h0;  // 32'h18e98ec8;
    ram_cell[     139] = 32'h0;  // 32'h9ae666da;
    ram_cell[     140] = 32'h0;  // 32'h94f6c982;
    ram_cell[     141] = 32'h0;  // 32'h0a2a0461;
    ram_cell[     142] = 32'h0;  // 32'h7ec90f88;
    ram_cell[     143] = 32'h0;  // 32'heef30d55;
    ram_cell[     144] = 32'h0;  // 32'hcf433698;
    ram_cell[     145] = 32'h0;  // 32'hfd90766d;
    ram_cell[     146] = 32'h0;  // 32'hdf40bf0b;
    ram_cell[     147] = 32'h0;  // 32'h0a40c41a;
    ram_cell[     148] = 32'h0;  // 32'h2651a747;
    ram_cell[     149] = 32'h0;  // 32'h3be0136e;
    ram_cell[     150] = 32'h0;  // 32'hcd10ce6c;
    ram_cell[     151] = 32'h0;  // 32'h921c55b3;
    ram_cell[     152] = 32'h0;  // 32'h437220b0;
    ram_cell[     153] = 32'h0;  // 32'he731d420;
    ram_cell[     154] = 32'h0;  // 32'h37d6f98c;
    ram_cell[     155] = 32'h0;  // 32'h8c7689c2;
    ram_cell[     156] = 32'h0;  // 32'h4084fcb7;
    ram_cell[     157] = 32'h0;  // 32'hbd970db6;
    ram_cell[     158] = 32'h0;  // 32'h9ae9d67d;
    ram_cell[     159] = 32'h0;  // 32'h10807ade;
    ram_cell[     160] = 32'h0;  // 32'h0b176dac;
    ram_cell[     161] = 32'h0;  // 32'ha30b119c;
    ram_cell[     162] = 32'h0;  // 32'hf4d97081;
    ram_cell[     163] = 32'h0;  // 32'hd8f8f890;
    ram_cell[     164] = 32'h0;  // 32'h658869d4;
    ram_cell[     165] = 32'h0;  // 32'h8a6d5714;
    ram_cell[     166] = 32'h0;  // 32'h6e9379af;
    ram_cell[     167] = 32'h0;  // 32'hfa9e086d;
    ram_cell[     168] = 32'h0;  // 32'h70116333;
    ram_cell[     169] = 32'h0;  // 32'hc8713823;
    ram_cell[     170] = 32'h0;  // 32'h5f754398;
    ram_cell[     171] = 32'h0;  // 32'hecc6c2a9;
    ram_cell[     172] = 32'h0;  // 32'h47ad46d2;
    ram_cell[     173] = 32'h0;  // 32'ha72bb86b;
    ram_cell[     174] = 32'h0;  // 32'h9b1b5019;
    ram_cell[     175] = 32'h0;  // 32'h15b84cc0;
    ram_cell[     176] = 32'h0;  // 32'h7cf474f8;
    ram_cell[     177] = 32'h0;  // 32'hce30f6c4;
    ram_cell[     178] = 32'h0;  // 32'h53869763;
    ram_cell[     179] = 32'h0;  // 32'h01a7d28d;
    ram_cell[     180] = 32'h0;  // 32'h2f8572f3;
    ram_cell[     181] = 32'h0;  // 32'h35112c88;
    ram_cell[     182] = 32'h0;  // 32'h650da12c;
    ram_cell[     183] = 32'h0;  // 32'hcffc37d0;
    ram_cell[     184] = 32'h0;  // 32'h00c3898a;
    ram_cell[     185] = 32'h0;  // 32'h9a9e5c65;
    ram_cell[     186] = 32'h0;  // 32'h7a734d7c;
    ram_cell[     187] = 32'h0;  // 32'h4e9cf466;
    ram_cell[     188] = 32'h0;  // 32'h76754c9c;
    ram_cell[     189] = 32'h0;  // 32'h619c06b3;
    ram_cell[     190] = 32'h0;  // 32'hae4049fe;
    ram_cell[     191] = 32'h0;  // 32'hce3f9f5e;
    ram_cell[     192] = 32'h0;  // 32'h51780c01;
    ram_cell[     193] = 32'h0;  // 32'hf40e4a90;
    ram_cell[     194] = 32'h0;  // 32'h28ddd62e;
    ram_cell[     195] = 32'h0;  // 32'hd31945e3;
    ram_cell[     196] = 32'h0;  // 32'h56153d58;
    ram_cell[     197] = 32'h0;  // 32'h570147cd;
    ram_cell[     198] = 32'h0;  // 32'h22c73cb2;
    ram_cell[     199] = 32'h0;  // 32'h035235a9;
    ram_cell[     200] = 32'h0;  // 32'hfafc8ed9;
    ram_cell[     201] = 32'h0;  // 32'h11721be9;
    ram_cell[     202] = 32'h0;  // 32'hd1d1005c;
    ram_cell[     203] = 32'h0;  // 32'hbd33ff66;
    ram_cell[     204] = 32'h0;  // 32'h5f68ab36;
    ram_cell[     205] = 32'h0;  // 32'h00855651;
    ram_cell[     206] = 32'h0;  // 32'hdc7da74d;
    ram_cell[     207] = 32'h0;  // 32'hb5ea9e20;
    ram_cell[     208] = 32'h0;  // 32'h5a62180f;
    ram_cell[     209] = 32'h0;  // 32'h4174f5d1;
    ram_cell[     210] = 32'h0;  // 32'h28c087b7;
    ram_cell[     211] = 32'h0;  // 32'h297c0ca9;
    ram_cell[     212] = 32'h0;  // 32'hdb918154;
    ram_cell[     213] = 32'h0;  // 32'hb7290dd5;
    ram_cell[     214] = 32'h0;  // 32'hc853fdcf;
    ram_cell[     215] = 32'h0;  // 32'hf27bd536;
    ram_cell[     216] = 32'h0;  // 32'hc336b70f;
    ram_cell[     217] = 32'h0;  // 32'ha55cc71c;
    ram_cell[     218] = 32'h0;  // 32'h74e10783;
    ram_cell[     219] = 32'h0;  // 32'he469596a;
    ram_cell[     220] = 32'h0;  // 32'hfdf02a12;
    ram_cell[     221] = 32'h0;  // 32'h24392f24;
    ram_cell[     222] = 32'h0;  // 32'hc44a8e90;
    ram_cell[     223] = 32'h0;  // 32'h6be7eedb;
    ram_cell[     224] = 32'h0;  // 32'h3e617473;
    ram_cell[     225] = 32'h0;  // 32'hf13ef30d;
    ram_cell[     226] = 32'h0;  // 32'hb1d89657;
    ram_cell[     227] = 32'h0;  // 32'he5604c7e;
    ram_cell[     228] = 32'h0;  // 32'h809982ad;
    ram_cell[     229] = 32'h0;  // 32'hc7327738;
    ram_cell[     230] = 32'h0;  // 32'hf95b3af6;
    ram_cell[     231] = 32'h0;  // 32'h1b242115;
    ram_cell[     232] = 32'h0;  // 32'hbcd12335;
    ram_cell[     233] = 32'h0;  // 32'h32374744;
    ram_cell[     234] = 32'h0;  // 32'h22cee06b;
    ram_cell[     235] = 32'h0;  // 32'h0cfd0625;
    ram_cell[     236] = 32'h0;  // 32'h39cc7eac;
    ram_cell[     237] = 32'h0;  // 32'hea606b9c;
    ram_cell[     238] = 32'h0;  // 32'hd9d7f68d;
    ram_cell[     239] = 32'h0;  // 32'ha5064c17;
    ram_cell[     240] = 32'h0;  // 32'hd8d9b4eb;
    ram_cell[     241] = 32'h0;  // 32'he6b17810;
    ram_cell[     242] = 32'h0;  // 32'h0dfc431d;
    ram_cell[     243] = 32'h0;  // 32'h4e207418;
    ram_cell[     244] = 32'h0;  // 32'h7fc07199;
    ram_cell[     245] = 32'h0;  // 32'h1eeadf79;
    ram_cell[     246] = 32'h0;  // 32'h25c8eea1;
    ram_cell[     247] = 32'h0;  // 32'h610250bf;
    ram_cell[     248] = 32'h0;  // 32'h55572db5;
    ram_cell[     249] = 32'h0;  // 32'h6c54f5be;
    ram_cell[     250] = 32'h0;  // 32'h94d7446d;
    ram_cell[     251] = 32'h0;  // 32'h969093e5;
    ram_cell[     252] = 32'h0;  // 32'hc7d9031a;
    ram_cell[     253] = 32'h0;  // 32'h856dc199;
    ram_cell[     254] = 32'h0;  // 32'hec139286;
    ram_cell[     255] = 32'h0;  // 32'h9179d667;
    // src matrix A
    ram_cell[     256] = 32'h916a52c2;
    ram_cell[     257] = 32'h8aa1f604;
    ram_cell[     258] = 32'hd13c1e22;
    ram_cell[     259] = 32'h28cfd377;
    ram_cell[     260] = 32'h5c17b23b;
    ram_cell[     261] = 32'hb3ff53a8;
    ram_cell[     262] = 32'h3c2b9291;
    ram_cell[     263] = 32'he69f79d3;
    ram_cell[     264] = 32'hf390219e;
    ram_cell[     265] = 32'h14327195;
    ram_cell[     266] = 32'h8ba0f8c2;
    ram_cell[     267] = 32'h1044acd0;
    ram_cell[     268] = 32'h0dd565c9;
    ram_cell[     269] = 32'hf905977a;
    ram_cell[     270] = 32'ha06d3870;
    ram_cell[     271] = 32'h38436ae1;
    ram_cell[     272] = 32'ha6376a56;
    ram_cell[     273] = 32'h45448147;
    ram_cell[     274] = 32'h94ddaa03;
    ram_cell[     275] = 32'hcec2ef0b;
    ram_cell[     276] = 32'h0b351f1a;
    ram_cell[     277] = 32'h6404884b;
    ram_cell[     278] = 32'h5d055509;
    ram_cell[     279] = 32'hc53278ec;
    ram_cell[     280] = 32'h819983a6;
    ram_cell[     281] = 32'h37ce720e;
    ram_cell[     282] = 32'hea7c3108;
    ram_cell[     283] = 32'hf9cd561f;
    ram_cell[     284] = 32'h09185396;
    ram_cell[     285] = 32'he6904911;
    ram_cell[     286] = 32'hbaf73107;
    ram_cell[     287] = 32'he3243b45;
    ram_cell[     288] = 32'h5286a4f1;
    ram_cell[     289] = 32'h37ba446e;
    ram_cell[     290] = 32'hb3b5cd7f;
    ram_cell[     291] = 32'h47fe5828;
    ram_cell[     292] = 32'h448e0a5f;
    ram_cell[     293] = 32'h6a64f4b4;
    ram_cell[     294] = 32'ha66f6a1d;
    ram_cell[     295] = 32'he96a3f5e;
    ram_cell[     296] = 32'h9c656745;
    ram_cell[     297] = 32'hb6589977;
    ram_cell[     298] = 32'hc1a0171d;
    ram_cell[     299] = 32'hbe1ca41b;
    ram_cell[     300] = 32'hc38ce590;
    ram_cell[     301] = 32'h164319b3;
    ram_cell[     302] = 32'h25deb749;
    ram_cell[     303] = 32'hc1e55e5d;
    ram_cell[     304] = 32'hd8aeec74;
    ram_cell[     305] = 32'h5c4e574e;
    ram_cell[     306] = 32'h2953dcef;
    ram_cell[     307] = 32'ha34ad383;
    ram_cell[     308] = 32'h73c96294;
    ram_cell[     309] = 32'h096d5d6d;
    ram_cell[     310] = 32'h6de2697d;
    ram_cell[     311] = 32'hc9af28b2;
    ram_cell[     312] = 32'h87a41d27;
    ram_cell[     313] = 32'hf8dfa4d9;
    ram_cell[     314] = 32'hefd72d36;
    ram_cell[     315] = 32'he4b446a9;
    ram_cell[     316] = 32'hd127c8b6;
    ram_cell[     317] = 32'habf01adf;
    ram_cell[     318] = 32'hf8e21ec6;
    ram_cell[     319] = 32'ha739481c;
    ram_cell[     320] = 32'h4333b645;
    ram_cell[     321] = 32'hceb82ce6;
    ram_cell[     322] = 32'h9e98eaef;
    ram_cell[     323] = 32'h9feadd7a;
    ram_cell[     324] = 32'h23013fe9;
    ram_cell[     325] = 32'hc7bfb7a5;
    ram_cell[     326] = 32'he5ff8f79;
    ram_cell[     327] = 32'he9df8225;
    ram_cell[     328] = 32'h475d3238;
    ram_cell[     329] = 32'h796f4b96;
    ram_cell[     330] = 32'hef5817e3;
    ram_cell[     331] = 32'h82064a38;
    ram_cell[     332] = 32'h12e7039f;
    ram_cell[     333] = 32'h84f39bb0;
    ram_cell[     334] = 32'h9011b750;
    ram_cell[     335] = 32'h73dd5540;
    ram_cell[     336] = 32'h9ae40a49;
    ram_cell[     337] = 32'h73ee2922;
    ram_cell[     338] = 32'h0ba42f22;
    ram_cell[     339] = 32'h679a6572;
    ram_cell[     340] = 32'h4b7655a5;
    ram_cell[     341] = 32'h33893cda;
    ram_cell[     342] = 32'h92aff5d5;
    ram_cell[     343] = 32'h1ba3276b;
    ram_cell[     344] = 32'h5102712e;
    ram_cell[     345] = 32'h68be7772;
    ram_cell[     346] = 32'h86cd0557;
    ram_cell[     347] = 32'hd622bca8;
    ram_cell[     348] = 32'h42e9a27d;
    ram_cell[     349] = 32'h1ce1ebbb;
    ram_cell[     350] = 32'h699db9f4;
    ram_cell[     351] = 32'hc5407080;
    ram_cell[     352] = 32'hccc3d9bd;
    ram_cell[     353] = 32'hb6c7e787;
    ram_cell[     354] = 32'h636a76e8;
    ram_cell[     355] = 32'h78906c0c;
    ram_cell[     356] = 32'h8cbd294d;
    ram_cell[     357] = 32'hf4dfd0c5;
    ram_cell[     358] = 32'hc769f367;
    ram_cell[     359] = 32'h1008386d;
    ram_cell[     360] = 32'h098224db;
    ram_cell[     361] = 32'h33a10c8c;
    ram_cell[     362] = 32'hcca4d923;
    ram_cell[     363] = 32'hbf36e373;
    ram_cell[     364] = 32'h56ce7e87;
    ram_cell[     365] = 32'hf49b8221;
    ram_cell[     366] = 32'h32499e2a;
    ram_cell[     367] = 32'h6b15e38f;
    ram_cell[     368] = 32'h40e619a7;
    ram_cell[     369] = 32'ha8d25aca;
    ram_cell[     370] = 32'hb4af8923;
    ram_cell[     371] = 32'hfea4d6a6;
    ram_cell[     372] = 32'h4bbabce2;
    ram_cell[     373] = 32'hed407db7;
    ram_cell[     374] = 32'h6fe44e47;
    ram_cell[     375] = 32'h494d615b;
    ram_cell[     376] = 32'ha8fdd3b3;
    ram_cell[     377] = 32'h2e6ee797;
    ram_cell[     378] = 32'hc63774a4;
    ram_cell[     379] = 32'hdcf240f0;
    ram_cell[     380] = 32'h6caf64ac;
    ram_cell[     381] = 32'h8c1b200d;
    ram_cell[     382] = 32'h918f8407;
    ram_cell[     383] = 32'h1103577a;
    ram_cell[     384] = 32'h9cbb94f7;
    ram_cell[     385] = 32'h24dbb03e;
    ram_cell[     386] = 32'h84b05c88;
    ram_cell[     387] = 32'h2aaf8e12;
    ram_cell[     388] = 32'hcfbba0db;
    ram_cell[     389] = 32'h246bf877;
    ram_cell[     390] = 32'h1b20f13d;
    ram_cell[     391] = 32'hf82a764b;
    ram_cell[     392] = 32'h97999fdf;
    ram_cell[     393] = 32'hca41aa53;
    ram_cell[     394] = 32'h3de9c445;
    ram_cell[     395] = 32'h913dcdb2;
    ram_cell[     396] = 32'h275d6784;
    ram_cell[     397] = 32'hfd901120;
    ram_cell[     398] = 32'h50a6564a;
    ram_cell[     399] = 32'h332b5066;
    ram_cell[     400] = 32'h27adec55;
    ram_cell[     401] = 32'h6053201b;
    ram_cell[     402] = 32'hfb7a60be;
    ram_cell[     403] = 32'ha90a6301;
    ram_cell[     404] = 32'hfbebb568;
    ram_cell[     405] = 32'h4112d42d;
    ram_cell[     406] = 32'h52765eb0;
    ram_cell[     407] = 32'h7eccb941;
    ram_cell[     408] = 32'h668dc785;
    ram_cell[     409] = 32'h6b2cd24f;
    ram_cell[     410] = 32'h94ca90e3;
    ram_cell[     411] = 32'h24ae25d1;
    ram_cell[     412] = 32'h4c42bf8d;
    ram_cell[     413] = 32'h25420485;
    ram_cell[     414] = 32'hd0512415;
    ram_cell[     415] = 32'h8a2be7f5;
    ram_cell[     416] = 32'hbdf8530c;
    ram_cell[     417] = 32'hb7b0cc09;
    ram_cell[     418] = 32'ha45b6b63;
    ram_cell[     419] = 32'h9b2d07b5;
    ram_cell[     420] = 32'h59b0f3dc;
    ram_cell[     421] = 32'hb91ff0ee;
    ram_cell[     422] = 32'hf563ac65;
    ram_cell[     423] = 32'h210587ac;
    ram_cell[     424] = 32'h006dad41;
    ram_cell[     425] = 32'h90a87f9b;
    ram_cell[     426] = 32'h826fc982;
    ram_cell[     427] = 32'h43161f0b;
    ram_cell[     428] = 32'h8f49d879;
    ram_cell[     429] = 32'hedf4392f;
    ram_cell[     430] = 32'h27d65cfd;
    ram_cell[     431] = 32'h7dc7f0bf;
    ram_cell[     432] = 32'ha0536e1f;
    ram_cell[     433] = 32'hb6fc07a8;
    ram_cell[     434] = 32'h4f993d17;
    ram_cell[     435] = 32'h5f3fd46c;
    ram_cell[     436] = 32'h12d290df;
    ram_cell[     437] = 32'hf2014f9a;
    ram_cell[     438] = 32'h5f85af1f;
    ram_cell[     439] = 32'h357e3052;
    ram_cell[     440] = 32'h7930b5b0;
    ram_cell[     441] = 32'h0fc76101;
    ram_cell[     442] = 32'h695d12df;
    ram_cell[     443] = 32'h474f1afd;
    ram_cell[     444] = 32'h1ebf2949;
    ram_cell[     445] = 32'h32f67246;
    ram_cell[     446] = 32'hd548e299;
    ram_cell[     447] = 32'he3ca6326;
    ram_cell[     448] = 32'h83b7aeab;
    ram_cell[     449] = 32'h6aef0ccf;
    ram_cell[     450] = 32'hdbc32267;
    ram_cell[     451] = 32'h53a8e7f7;
    ram_cell[     452] = 32'h1496e0ff;
    ram_cell[     453] = 32'hefb2f9da;
    ram_cell[     454] = 32'h74503dc2;
    ram_cell[     455] = 32'hccf9ab46;
    ram_cell[     456] = 32'h4f6d3fba;
    ram_cell[     457] = 32'h959e30ed;
    ram_cell[     458] = 32'h3a1b1e06;
    ram_cell[     459] = 32'h55340aa2;
    ram_cell[     460] = 32'he1167c67;
    ram_cell[     461] = 32'hac10cd32;
    ram_cell[     462] = 32'h821faaf7;
    ram_cell[     463] = 32'h4003ac18;
    ram_cell[     464] = 32'h898db45d;
    ram_cell[     465] = 32'h3f884631;
    ram_cell[     466] = 32'h26786677;
    ram_cell[     467] = 32'h6d2eee88;
    ram_cell[     468] = 32'h15924894;
    ram_cell[     469] = 32'h4c0b55a4;
    ram_cell[     470] = 32'h65e35fc8;
    ram_cell[     471] = 32'haf334724;
    ram_cell[     472] = 32'hbba06fa5;
    ram_cell[     473] = 32'h2529675a;
    ram_cell[     474] = 32'h2c1a51d3;
    ram_cell[     475] = 32'hb78eb297;
    ram_cell[     476] = 32'h989efb5e;
    ram_cell[     477] = 32'h978eb7f5;
    ram_cell[     478] = 32'h4da9cca6;
    ram_cell[     479] = 32'hd3002fa7;
    ram_cell[     480] = 32'hf21b6da6;
    ram_cell[     481] = 32'h3a4fc718;
    ram_cell[     482] = 32'h3f5e8ba4;
    ram_cell[     483] = 32'hf0e240d4;
    ram_cell[     484] = 32'h41217176;
    ram_cell[     485] = 32'h82884c45;
    ram_cell[     486] = 32'hc88332ba;
    ram_cell[     487] = 32'h15fc3546;
    ram_cell[     488] = 32'h67f2790c;
    ram_cell[     489] = 32'hc4a749d3;
    ram_cell[     490] = 32'h5faea486;
    ram_cell[     491] = 32'he72038a0;
    ram_cell[     492] = 32'hc3c4cb6d;
    ram_cell[     493] = 32'he1d64507;
    ram_cell[     494] = 32'hdf2413f3;
    ram_cell[     495] = 32'h0af70863;
    ram_cell[     496] = 32'hb4a06da5;
    ram_cell[     497] = 32'h7f61f6a9;
    ram_cell[     498] = 32'h7a528525;
    ram_cell[     499] = 32'h397e2d9d;
    ram_cell[     500] = 32'hc4038c2d;
    ram_cell[     501] = 32'hdf7a496c;
    ram_cell[     502] = 32'h326f0627;
    ram_cell[     503] = 32'hd4647d9c;
    ram_cell[     504] = 32'hd626812f;
    ram_cell[     505] = 32'h7d53024a;
    ram_cell[     506] = 32'hf41f5f63;
    ram_cell[     507] = 32'h2c03b8c6;
    ram_cell[     508] = 32'h60f30414;
    ram_cell[     509] = 32'h991e0cff;
    ram_cell[     510] = 32'hc599a056;
    ram_cell[     511] = 32'h12ed313f;
    // src matrix B
    ram_cell[     512] = 32'h310a1f01;
    ram_cell[     513] = 32'hfe7806eb;
    ram_cell[     514] = 32'hb50aa23d;
    ram_cell[     515] = 32'h0bc9852e;
    ram_cell[     516] = 32'hbd2f88d8;
    ram_cell[     517] = 32'hb9645ad2;
    ram_cell[     518] = 32'had9fb53f;
    ram_cell[     519] = 32'h5bd9f27a;
    ram_cell[     520] = 32'h014a6f5b;
    ram_cell[     521] = 32'hddc38444;
    ram_cell[     522] = 32'hac9596f0;
    ram_cell[     523] = 32'h4fb7a5fc;
    ram_cell[     524] = 32'hf198a123;
    ram_cell[     525] = 32'ha2c7c785;
    ram_cell[     526] = 32'hc596a8b8;
    ram_cell[     527] = 32'h772f2cec;
    ram_cell[     528] = 32'h312b7b73;
    ram_cell[     529] = 32'hfd050944;
    ram_cell[     530] = 32'h367ee0fa;
    ram_cell[     531] = 32'hf09422d5;
    ram_cell[     532] = 32'h064021c4;
    ram_cell[     533] = 32'h50a62510;
    ram_cell[     534] = 32'h7d253e47;
    ram_cell[     535] = 32'h7ce47f2d;
    ram_cell[     536] = 32'h3ca5b302;
    ram_cell[     537] = 32'h7e3efb99;
    ram_cell[     538] = 32'h692eadde;
    ram_cell[     539] = 32'h92f79195;
    ram_cell[     540] = 32'h76156b0a;
    ram_cell[     541] = 32'hddebb72b;
    ram_cell[     542] = 32'h2ab9fdc2;
    ram_cell[     543] = 32'h43cb3f21;
    ram_cell[     544] = 32'h9051d396;
    ram_cell[     545] = 32'h9f9c8d33;
    ram_cell[     546] = 32'hcbe2723f;
    ram_cell[     547] = 32'hc679c7cc;
    ram_cell[     548] = 32'hca71b8c0;
    ram_cell[     549] = 32'h1fd3d5d3;
    ram_cell[     550] = 32'he71a23db;
    ram_cell[     551] = 32'hc33df237;
    ram_cell[     552] = 32'h64d0430b;
    ram_cell[     553] = 32'h5438af7b;
    ram_cell[     554] = 32'h4f409b90;
    ram_cell[     555] = 32'h2f4490f0;
    ram_cell[     556] = 32'h8e3ae29d;
    ram_cell[     557] = 32'h89f92876;
    ram_cell[     558] = 32'h6a72a826;
    ram_cell[     559] = 32'h72fb93c7;
    ram_cell[     560] = 32'ha7dc94b1;
    ram_cell[     561] = 32'h61657a71;
    ram_cell[     562] = 32'he541751e;
    ram_cell[     563] = 32'hf01a5ddf;
    ram_cell[     564] = 32'hf01406f9;
    ram_cell[     565] = 32'he0f45b54;
    ram_cell[     566] = 32'h5874154e;
    ram_cell[     567] = 32'h69208997;
    ram_cell[     568] = 32'h74402ed9;
    ram_cell[     569] = 32'hd21b8432;
    ram_cell[     570] = 32'h4bb214d9;
    ram_cell[     571] = 32'h848de975;
    ram_cell[     572] = 32'h90583b3f;
    ram_cell[     573] = 32'h81c403b9;
    ram_cell[     574] = 32'h00b2a3bd;
    ram_cell[     575] = 32'hfe5d61c3;
    ram_cell[     576] = 32'hae12336e;
    ram_cell[     577] = 32'h88bf8b34;
    ram_cell[     578] = 32'h06692853;
    ram_cell[     579] = 32'hac2aff2c;
    ram_cell[     580] = 32'h092933a9;
    ram_cell[     581] = 32'h7b6d369a;
    ram_cell[     582] = 32'h2a4ef82c;
    ram_cell[     583] = 32'h12a942ea;
    ram_cell[     584] = 32'h49cff434;
    ram_cell[     585] = 32'hcdf1d778;
    ram_cell[     586] = 32'hf6e7785c;
    ram_cell[     587] = 32'h30a22b82;
    ram_cell[     588] = 32'h90344ce8;
    ram_cell[     589] = 32'hbbfd9b75;
    ram_cell[     590] = 32'h67c04d92;
    ram_cell[     591] = 32'h6557d4cf;
    ram_cell[     592] = 32'h557de6d5;
    ram_cell[     593] = 32'h4be45223;
    ram_cell[     594] = 32'hadd422fd;
    ram_cell[     595] = 32'h15bf8556;
    ram_cell[     596] = 32'hc36cd058;
    ram_cell[     597] = 32'h58393814;
    ram_cell[     598] = 32'hd01153cc;
    ram_cell[     599] = 32'h96135946;
    ram_cell[     600] = 32'h4493b093;
    ram_cell[     601] = 32'h67b80217;
    ram_cell[     602] = 32'hbe137989;
    ram_cell[     603] = 32'he6eee272;
    ram_cell[     604] = 32'hce421e4f;
    ram_cell[     605] = 32'h0c236f9b;
    ram_cell[     606] = 32'had0c44dd;
    ram_cell[     607] = 32'h5cb5f120;
    ram_cell[     608] = 32'heaa14b15;
    ram_cell[     609] = 32'hb4553219;
    ram_cell[     610] = 32'h714c7ed4;
    ram_cell[     611] = 32'h758ccb99;
    ram_cell[     612] = 32'hbd91dada;
    ram_cell[     613] = 32'h6623e858;
    ram_cell[     614] = 32'ha5a37ebf;
    ram_cell[     615] = 32'hddadd90d;
    ram_cell[     616] = 32'h03c19717;
    ram_cell[     617] = 32'h115fc917;
    ram_cell[     618] = 32'hac6d77b1;
    ram_cell[     619] = 32'h041f421e;
    ram_cell[     620] = 32'hb3768c5f;
    ram_cell[     621] = 32'h531ccae7;
    ram_cell[     622] = 32'h68fe3699;
    ram_cell[     623] = 32'hf9cdbe34;
    ram_cell[     624] = 32'hcf0c7bc9;
    ram_cell[     625] = 32'h34d4c42a;
    ram_cell[     626] = 32'hc0ee20c5;
    ram_cell[     627] = 32'h649217bb;
    ram_cell[     628] = 32'h05996474;
    ram_cell[     629] = 32'h4d253c44;
    ram_cell[     630] = 32'h288fa86d;
    ram_cell[     631] = 32'h06d1726b;
    ram_cell[     632] = 32'hed52ca18;
    ram_cell[     633] = 32'h4186827d;
    ram_cell[     634] = 32'hefefd5e6;
    ram_cell[     635] = 32'h226ef525;
    ram_cell[     636] = 32'h4650b631;
    ram_cell[     637] = 32'h4dbd59f5;
    ram_cell[     638] = 32'he4fee7bf;
    ram_cell[     639] = 32'h565c7d27;
    ram_cell[     640] = 32'heecea009;
    ram_cell[     641] = 32'hfc1dc718;
    ram_cell[     642] = 32'hdafb6599;
    ram_cell[     643] = 32'h5dbc35b6;
    ram_cell[     644] = 32'ha1207aa1;
    ram_cell[     645] = 32'hb99ae13f;
    ram_cell[     646] = 32'hfb680b3b;
    ram_cell[     647] = 32'hf7646063;
    ram_cell[     648] = 32'hc4b644a0;
    ram_cell[     649] = 32'h37c309ec;
    ram_cell[     650] = 32'h5cfbe1ca;
    ram_cell[     651] = 32'h3855b77a;
    ram_cell[     652] = 32'h2dad88b6;
    ram_cell[     653] = 32'hf37b523d;
    ram_cell[     654] = 32'hc41f59a1;
    ram_cell[     655] = 32'h824e0e22;
    ram_cell[     656] = 32'h48d727d5;
    ram_cell[     657] = 32'hc8b13298;
    ram_cell[     658] = 32'h0a3cb787;
    ram_cell[     659] = 32'hd5147bb2;
    ram_cell[     660] = 32'h0535ce86;
    ram_cell[     661] = 32'h6b7b9ab3;
    ram_cell[     662] = 32'h7996eccc;
    ram_cell[     663] = 32'h4394a237;
    ram_cell[     664] = 32'h9da14c34;
    ram_cell[     665] = 32'h34518a57;
    ram_cell[     666] = 32'h4d8c038e;
    ram_cell[     667] = 32'h01a8a821;
    ram_cell[     668] = 32'h26f172c4;
    ram_cell[     669] = 32'h6486fcc8;
    ram_cell[     670] = 32'hfd2ae763;
    ram_cell[     671] = 32'h3e7903e9;
    ram_cell[     672] = 32'hc41c1584;
    ram_cell[     673] = 32'h7e6597b5;
    ram_cell[     674] = 32'h5cc7a516;
    ram_cell[     675] = 32'h8cc13012;
    ram_cell[     676] = 32'hcfc761f5;
    ram_cell[     677] = 32'had94550b;
    ram_cell[     678] = 32'h4e09ef99;
    ram_cell[     679] = 32'h190b7b7b;
    ram_cell[     680] = 32'h39e0c5d5;
    ram_cell[     681] = 32'h041cb13d;
    ram_cell[     682] = 32'h9b96141c;
    ram_cell[     683] = 32'h52ece100;
    ram_cell[     684] = 32'hc23b39ea;
    ram_cell[     685] = 32'hfc7215c9;
    ram_cell[     686] = 32'h1b9ea649;
    ram_cell[     687] = 32'hec3de9a2;
    ram_cell[     688] = 32'hb331fd14;
    ram_cell[     689] = 32'h3cafd7b9;
    ram_cell[     690] = 32'h51756a13;
    ram_cell[     691] = 32'ha7e53d93;
    ram_cell[     692] = 32'he1f6d575;
    ram_cell[     693] = 32'h792a9462;
    ram_cell[     694] = 32'hf88c3aeb;
    ram_cell[     695] = 32'hc39d204f;
    ram_cell[     696] = 32'hb1bafd1e;
    ram_cell[     697] = 32'hc29872c7;
    ram_cell[     698] = 32'hb46e99c6;
    ram_cell[     699] = 32'h4df78cdc;
    ram_cell[     700] = 32'hf5d32a98;
    ram_cell[     701] = 32'hfa3aa858;
    ram_cell[     702] = 32'hd3e00974;
    ram_cell[     703] = 32'h0770df8c;
    ram_cell[     704] = 32'h0bceb430;
    ram_cell[     705] = 32'h7b89b009;
    ram_cell[     706] = 32'h542fbb62;
    ram_cell[     707] = 32'h9fb3f451;
    ram_cell[     708] = 32'hc9144ae4;
    ram_cell[     709] = 32'hd1b45778;
    ram_cell[     710] = 32'h0a9bf478;
    ram_cell[     711] = 32'hcf7b8196;
    ram_cell[     712] = 32'h5cf01ce6;
    ram_cell[     713] = 32'h2b4f955b;
    ram_cell[     714] = 32'h8c76678b;
    ram_cell[     715] = 32'hcafa3a42;
    ram_cell[     716] = 32'hbe5b56fd;
    ram_cell[     717] = 32'h1c5f3e1e;
    ram_cell[     718] = 32'h52de3c58;
    ram_cell[     719] = 32'h18d35caa;
    ram_cell[     720] = 32'hc6ce82c4;
    ram_cell[     721] = 32'hefface1c;
    ram_cell[     722] = 32'ha317cfc3;
    ram_cell[     723] = 32'ha98ee5e9;
    ram_cell[     724] = 32'hb93caa33;
    ram_cell[     725] = 32'haf1a2204;
    ram_cell[     726] = 32'h13d90805;
    ram_cell[     727] = 32'h42f8ab1e;
    ram_cell[     728] = 32'h8c89de1a;
    ram_cell[     729] = 32'h18924a38;
    ram_cell[     730] = 32'h66f7b6e0;
    ram_cell[     731] = 32'hcd2ba8c1;
    ram_cell[     732] = 32'h94a9f15b;
    ram_cell[     733] = 32'h230f6605;
    ram_cell[     734] = 32'h8a14463a;
    ram_cell[     735] = 32'h120de06c;
    ram_cell[     736] = 32'h0ac2d497;
    ram_cell[     737] = 32'hf98b9d88;
    ram_cell[     738] = 32'h5e5ea146;
    ram_cell[     739] = 32'h8a4bff92;
    ram_cell[     740] = 32'h228f6ffe;
    ram_cell[     741] = 32'h4dc67e17;
    ram_cell[     742] = 32'hd25854fd;
    ram_cell[     743] = 32'h74dc87eb;
    ram_cell[     744] = 32'h59e453e6;
    ram_cell[     745] = 32'h2716c40d;
    ram_cell[     746] = 32'ha6952fac;
    ram_cell[     747] = 32'h674f3e55;
    ram_cell[     748] = 32'h1ef3a5d2;
    ram_cell[     749] = 32'h5586f983;
    ram_cell[     750] = 32'h0ab91875;
    ram_cell[     751] = 32'h8b0ab9c9;
    ram_cell[     752] = 32'hd6a6e8c0;
    ram_cell[     753] = 32'haaee8563;
    ram_cell[     754] = 32'h829c5742;
    ram_cell[     755] = 32'h0feca812;
    ram_cell[     756] = 32'h39b32f24;
    ram_cell[     757] = 32'h70bdd8b4;
    ram_cell[     758] = 32'h1179cce4;
    ram_cell[     759] = 32'hf61cbb41;
    ram_cell[     760] = 32'hef6e0d4c;
    ram_cell[     761] = 32'h5638e410;
    ram_cell[     762] = 32'h1b8bd6f5;
    ram_cell[     763] = 32'h924bcd1e;
    ram_cell[     764] = 32'ha496a5bb;
    ram_cell[     765] = 32'h079b37b5;
    ram_cell[     766] = 32'h076d0536;
    ram_cell[     767] = 32'h3b4a468b;
end

endmodule